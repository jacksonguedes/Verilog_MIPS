module Desafio_ULA(input [3:0] a, b, input [1:0] selecao,
                   output reg [3:0] saida);
		always@(*)
			
			if (selecao == 2'b00)
				saida = a + b;
			else if (selecao == 2'b01)
				saida = a - b;
			else if (selecao == 2'b10)
				saida = a >> b;
			else if (selecao == 2'b11)
				saida = a << b;
	
endmodule
